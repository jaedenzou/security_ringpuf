`timescale 1ns / 1ps

//Comment out the line below while implementing your design with hard macro
(*KEEP_HIERARCHY="TRUE"*)

module ringoscillator(enable, reset, dffout);
    input enable, reset;
    output dffout;
	 
   //Comment out the line below while implementing your design with hard macro
	(* S = "TRUE" *)
	
	//Write the code for your ring oscillator
	//Comment it out after you create the hard macro



	/////////////////////////////////////////
	
endmodule